`ifndef AXI_SEQUENCER_SV
`define AXI_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer#(axi_tx) axi_sequencer_t;


`endif  // AXI_SEQUENCER_SV
